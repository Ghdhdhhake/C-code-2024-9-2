LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY count60 IS --60进制计数器
	PORT (
   		 CLK,RST,EN:IN STD_LOGIC;
   		 DHOUT:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0); --高四位输出
    	    DLOUT:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0); --低四位输出
         COUT:OUT STD_LOGIC);
END ENTITY count60;
ARCHITECTURE behave OF count60 IS
BEGIN
   COUT<='1'WHEN(DHOUT="0101" AND DLOUT="1001")ELSE '0'; --确定进位条件
	PROCESS(CLK,EN,RST)
	BEGIN
	      IF RST='1' THEN DHOUT<="0000";DLOUT<="0000"; --异步清零
	      ELSIF CLK'EVENT AND CLK ='1' THEN 
			IF EN='1' THEN DLOUT<=DLOUT+1;END IF;   --同步使能
			IF(DLOUT=9)THEN DLOUT<="0000";DHOUT<=DHOUT+1;END IF;  --低四位归零设置
	       IF(DHOUT=5 AND DLOUT=9) THEN DHOUT<="0000"; END IF; --高四位归零设置
			  END IF;
END PROCESS;
END ARCHITECTURE behave;