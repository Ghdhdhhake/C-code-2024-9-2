LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL ;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY smg IS  
	PORT (INDATA: IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		  ODATA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END ENTITY smg;
ARCHITECTURE BHV OF smg IS
	BEGIN
	PROCESS (INDATA)
	BEGIN
		CASE (INDATA) IS
			WHEN "0000" => ODATA<= "1000000" ; 
			WHEN "0001" => ODATA<= "1111001" ; 
			WHEN "0010" => ODATA<= "0100100" ; 
			WHEN "0011" => ODATA<= "0110000" ; 
			WHEN "0100" => ODATA<= "0011001" ; 
			WHEN "0101" => ODATA<= "0010010" ; 
			WHEN "0110" => ODATA<= "0000010" ; 
			WHEN "0111" => ODATA<= "1111000" ; 
			WHEN "1000" => ODATA<= "0000000" ; 
			WHEN "1001" => ODATA<= "0010000" ; 
			WHEN OTHERS => NULL;  
		END CASE; 
	END PROCESS;
END ARCHITECTURE BHV;